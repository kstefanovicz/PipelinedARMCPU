module flagReg(

  input logic


);
